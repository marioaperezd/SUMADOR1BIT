module C_XOR (A,B,OUT);
  input A,B;
  output OUT;
  
  assign OUT=A ^ B;
endmodule
