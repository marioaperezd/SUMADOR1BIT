module C_AND (A,B,OUT);
  input A,B;
  output OUT;
  
  assign OUT=A & B;
endmodule
